module explicit_types(
    input logic clk,
    input wire rst_n,
    output reg data_valid,
    inout tri data_bus
);
endmodule