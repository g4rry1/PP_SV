module vector_ports(
    input [7:0] data_bus,
    output [15:0] address_bus,
    inout [3:0] control_bus
);
endmodule