module signed_ports(
    input signed [15:0] signed_input,
    output signed [31:0] signed_output
);
endmodule