module no_parameters(input logic clk);
endmodule