module parent_module;
    child_module inst1(clk, rst, data_in, data_out);
endmodule