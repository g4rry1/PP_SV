module packed_arrays(
    input logic [3:0][7:0] packed_input,  // 4x8 бит
    output bit [2:0][15:0] packed_output  // 3x16 бит
);
endmodule