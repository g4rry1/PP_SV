module mixed_types(
    input logic a,      // logic input
    output wire b,      // wire output
    inout triand c      // triand inout
);
endmodule