(* optimize_power = "yes" *)
module attributed_module(
    input logic clk
);
endmodule