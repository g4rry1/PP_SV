module no_ports;
    logic internal_signal;
endmodule