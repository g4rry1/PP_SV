module interface_module(
    virtual bus_if bus_interface
);
endmodule