module single_bit(
    input bit a,
    output bit b
);
endmodule