module interface_instance(
    input clock_if clk_intf,
    output data_if data_intf
);
endmodule