module non_ansi_style(a, b, c);
    input a;
    output b;
    inout c;
    wire a, c;
    reg b;
endmodule