module implicit_types(
    input a,        // wire a
    output b,       // wire b
    inout c         // wire c
);
endmodule