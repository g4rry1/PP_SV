module with_parameters #(
    parameter WIDTH = 8,
    parameter DEPTH = 16
) (
    input logic [WIDTH-1:0] data_in,
    output logic [WIDTH-1:0] data_out
);
endmodule