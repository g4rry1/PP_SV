module parameterized_vectors #(
    parameter DATA_WIDTH = 32,
    parameter ADDR_WIDTH = 16
) (
    input [DATA_WIDTH-1:0] data_in,
    output [ADDR_WIDTH-1:0] addr_out
);
endmodule