module unpacked_arrays(
    input logic [7:0] array_input [0:3],  // 4 элемента по 8 бит
    output int array_output [8]           // 8 элементов по 32 бита
);
endmodule