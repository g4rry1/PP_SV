module value_parameters #(
    parameter WIDTH = 8,
    parameter real FREQUENCY = 100.0e6,
    parameter string MODULE_NAME = "default"
) (
    input [WIDTH-1:0] a
);
endmodule