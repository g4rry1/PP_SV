module top_level;
    sub_module inst1();
    another_module inst2();
endmodule

module sub_module;
    // содержимое
endmodule

module another_module;
    // содержимое
endmodule