module ansi_style(
    input a,
    output b,
    inout c
);
    // содержимое
endmodule